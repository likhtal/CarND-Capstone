camera_info:
  image_width: 800
  image_height: 600
stop_line_positions:
    - [1148.56, 1184.65]
    - [1559.2, 1158.43]
    - [2122.14, 1526.79]
    - [2175.237, 1795.71]
    - [1493.29, 2947.67]
    - [821.96, 2905.8]
    - [161.76, 2303.82]
    - [351.84, 1574.65]
manual_light_positions:
    - [1172.183, 1186.299, 5.576891]
    - [1584.065, 1156.953, 5.576705]
    - [2126.353, 1550.636, 5.576704]
    - [2178.291, 1819.328, 5.576704]
    - [1469.499, 2946.970, 5.576707]
    - [797.9147, 2905.590, 5.576708]
    - [160.8088, 2279.929, 5.606704]
    - [363.3780, 1553.731, 5.606708]